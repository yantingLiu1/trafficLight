library ieee;
use ieee.std_logic_1164.all;

entity synchronizer is
  port (
    clk   : in std_logic;
    reset : in std_logic;
    din   : in std_logic;
    dout  : out std_logic
  );
end synchronizer;

architecture circuit of synchronizer is
  signal sreg : std_logic_vector(1 downto 0);
begin

  sync_proc: process(clk, reset)
  begin
    if reset = '1' then
      sreg <= (others => '0');
    elsif rising_edge(clk) then
      sreg(0) <= din;
      sreg(1) <= sreg(0);
    end if;
  end process sync_proc;

  dout <= sreg(1);

end circuit;